// File Name: 32_MDR.v
`timescale 1ns/10ps
module Decoder4to16(
	input [3:0] decoderIn,
	output reg d0, d1, d2, d3, d4, d5, d6, d7, d8, d9, d10, d11, d12, d13, d14, d15);
	
	always @(decoderIn) begin
		case(decoderIn)
			4'b0000: begin 
				d0=1; d1=0; d2=0; d3=0; d4=0; d5=0; d6=0; d7=0; d8=0; d9=0; d10=0; d11=0; d12=0; d13=0; d14=0; d15=0; end

			4'b0001: begin 
				d0=0; d1=1; d2=0; d3=0; d4=0; d5=0; d6=0; d7=0; d8=0; d9=0; d10=0; d11=0; d12=0; d13=0; d14=0; d15=0; end
				
			4'b0010: begin d2=1; 
				d0=0; d1=0; d3=0; d4=0; d5=0; d6=0; d7=0; d8=0; d9=0; d10=0; d11=0; d12=0; d13=0; d14=0; d15=0; end
				
			4'b0011: begin d3=1; 
				d0=0; d1=0; d2=0; d4=0; d5=0; d6=0; d7=0; d8=0; d9=0; d10=0; d11=0; d12=0; d13=0; d14=0; d15=0; end
				
			4'b0100: begin d4=1; 
				d0=0; d1=0; d2=0; d3=0; d5=0; d6=0; d7=0; d8=0; d9=0; d10=0; d11=0; d12=0; d13=0; d14=0; d15=0; end
				
			4'b0101: begin d5=1; 
				d0=0; d1=0; d2=0; d3=0; d4=0;d6=0; d7=0; d8=0; d9=0; d10=0; d11=0; d12=0; d13=0; d14=0; d15=0; end
				
			4'b0110: begin d6=1; 
				d0=0; d1=0; d2=0; d3=0; d4=0; d5=0; d7=0; d8=0; d9=0; d10=0; d11=0; d12=0; d13=0; d14=0; d15=0; end
				
			4'b0111: begin d7=1; 
				d0=0; d1=0; d2=0; d3=0; d4=0; d5=0; d6=0;d8=0; d9=0; d10=0; d11=0; d12=0; d13=0; d14=0; d15=0; end
				
			4'b1000: begin d8=1; 
				d0=0; d1=0; d2=0; d3=0; d4=0; d5=0; d6=0; d7=0; d9=0; d10=0; d11=0; d12=0; d13=0; d14=0; d15=0; end
				
			4'b1001: begin d9=1; 
				d0=0; d1=0; d2=0; d3=0; d4=0; d5=0; d6=0; d7=0; d8=0; d10=0; d11=0; d12=0; d13=0; d14=0; d15=0; end
				
			4'b1010: begin d10=1; 
				d0=0; d1=0; d2=0; d3=0; d4=0; d5=0; d6=0; d7=0; d8=0; d9=0; d11=0; d12=0; d13=0; d14=0; d15=0; end
				
			4'b1011: begin d11=1; 
				d0=0; d1=0; d2=0; d3=0; d4=0; d5=0; d6=0; d7=0; d8=0; d9=0; d10=0; d12=0; d13=0; d14=0; d15=0; end
				
			4'b1100: begin d12=1; 
				d0=0; d1=0; d2=0; d3=0; d4=0; d5=0; d6=0; d7=0; d8=0; d9=0; d10=0; d11=0; d13=0; d14=0; d15=0; end
				
			4'b1101: begin d13=1; 
				d0=0; d1=0; d2=0; d3=0; d4=0; d5=0; d6=0; d7=0; d8=0; d9=0; d10=0; d11=0; d12=0; d14=0; d15=0; end
				
			4'b1110: begin d14=1; 
				d0=0; d1=0; d2=0; d3=0; d4=0; d5=0; d6=0; d7=0; d8=0; d9=0; d10=0; d11=0; d12=0; d13=0; d15=0; end
				
			4'b1111: begin d15=1; 
				d0=0; d1=0; d2=0; d3=0; d4=0; d5=0; d6=0; d7=0; d8=0; d9=0; d10=0; d11=0; d12=0; d13=0; d14=0; end
				
		endcase
	end
		
endmodule
